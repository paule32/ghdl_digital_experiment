------------------------------------------------------------------------------
-- File:    or_gate_7432.vhdl
-- Author:  (c) 2023 Jens Kallup - paule32
--
-- License: MIT - only for education, and non-profit !
------------------------------------------------------------------------------
-- used format:
-- ============
-- E_n => Eingang/Input  (Bsp: E_0, E_1, ...)
-- A_n => Ausgang/Output (Bsp: A_0 )
------------------------------------------------------------------------------
library ieee;

use ieee.std_logic_1164.all;
use work.Eingang2_Ausgang1_Record.all;

------------------------------------------------------------------------------
-- 7432 Quad 2-Eingangs-Logik ODER Gatter:
-- =======================================
--  Vcc
--    14 13 12     11   10  9      8
--     |  |  |      |    |  |      |
--     |  +  +      +    +  +      +
-- )---o--|--|------|----|--|------|---(
-- |      +  +      +    +  +      +   |
-- |      |  |      |    |  |      |   |
-- |      |  +--\   |    |  +--\   |   |
-- |      |      +--+    |      +--+   |
--  )     +-----/        +-----/       |
--  )                                  |
--  )  +-----\        +-----\          |
-- |   |      +--+    |      +--+      |
-- |   |  +--/   |    |  +--/   |      |
-- |   |  |      |    |  |      |      |
-- |   +  +      +    +  +      +      |
-- )---|--|------|----|--|------|--o---(
--     +  +      +    +  +      +  |
--     |  |      |    |  |      |  |
--     1  2      3    4  5      6  7 
--                                 Gnd
------------------------------------------------------------------------------
-- B => Block
-- A => Ausgang Port
-- E => Eingang Port
--
-- TTL ODER Gate:
-- ==============
-- B      1              2              3              4
-- A      3              6              8              11
-- E  1       2      4       5      9       10     12      13
------------------------------------------------------------------------------
--   E_0     E_1    E_2     E_3    E_4     E_5    E_6     E_7      E_0  +  E_1
--  ----- | -----  ----- | -----  ----- | -----  ----- | -----    ------------
--    0   |   0      0   |   0      0   |   0      0   |   0            0
--    0   |   1      0   |   1      0   |   1      0   |   1            1
--    1   |   0      1   |   0      1   |   0      1   |   0            1
--    1   |   1      1   |   1      1   |   1      1   |   1            1
------------------------------------------------------------------------------

------------------------------------------------------------------------------
-- Port-Zuweisung:
------------------------------------------------------------------------------
entity or_gate_7432 is
    port (
        Block_0 : in work.Eingang2_Ausgang1_Record.Bauteil;
        Block_1 : in work.Eingang2_Ausgang1_Record.Bauteil;
        Block_2 : in work.Eingang2_Ausgang1_Record.Bauteil;
        Block_3 : in work.Eingang2_Ausgang1_Record.Bauteil
    );
end entity or_gate_7432;

------------------------------------------------------------------------------
-- Architektur: Logik, und Signal-Verarbeitung
------------------------------------------------------------------------------
architecture or_7432_arch of or_gate_7432 is
begin
    process (Block_0, Block_1, Block_2, Block_3)
    begin
        Block_0.A_0 <= Block_0.E_0 or Block_0.E_1;
        Block_1.A_0 <= Block_1.E_0 or Block_1.E_1;
        Block_2.A_0 <= Block_2.E_0 or Block_2.E_1;
        Block_3.A_0 <= Block_3.E_0 or Block_3.E_1;
    end process;
end architecture or_7432_arch;

configuration or_7432_config of or_gate_7432 is
    for or_7432_arch
    end for;
end configuration or_7432_config;

------------------------------------------------------------------------------
-- E O F  -  End Of File.
------------------------------------------------------------------------------
