
library ieee;
use ieee.std_logic_1164.all;

package Eingang2_Ausgang1_Record is
    type Bauteil is record
        E_0 : std_logic;
        E_1 : std_logic;
        A_0 : std_logic;
    end record;
end package Eingang2_Ausgang1_Record;

-- Implementrierung
package body Eingang2_Ausgang1_Record is
end package body Eingang2_Ausgang1_Record;
